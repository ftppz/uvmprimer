/*
   Copyright 2013 Ray Salemi

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
*/
package example_pkg;
	import uvm_pkg::*;
`include "uvm_macros.svh"

	virtual clk_bfm clk_bfm_i;

`include "producer.svh"
`include "consumer.svh"
`include "communication_test.svh"
endpackage : example_pkg

   
     
   